
module register_file(input logic clk, rst, regWrite, 
							input logic [3:0] A1, A2, A3, 
							input logic [15:0] WD3, R15,
							output logic [15:0] RD1, RD2);
		// # bits         // # registros			
	logic [15:0] registers [15:0];
	logic [15:0] RD1_temp = 16'h0;
	logic [15:0] RD2_temp = 16'h0;
	
	
	// escritura se hace en flanco positivo
	always_ff @(posedge clk or posedge rst) begin
	
		if (rst) begin
			// Reset behavior
			registers[0] <= 16'd0;
			registers[1] <= 16'd0;
			registers[2] <= 16'd0;
			registers[3] <= 16'd0;
			registers[4] <= 16'd0;
			registers[5] <= 16'd0;
			registers[6] <= 16'd0;
			registers[7] <= 16'd0;
			registers[8] <= 16'd0;
			registers[9] <= 16'd0;
			registers[10] <= 16'd0;
			registers[11] <= 16'd0;
			registers[12] <= 16'd0; // registro de ubicación de pixeles (PU) 
			registers[13] <= 16'd0; // registro para la memoria (SP)
			registers[14] <= 16'd0; // registro para el contador del programa (PC)
			registers[15] <= 16'd0; //
		end 
		else begin
		
			if (regWrite) begin // si esta la senal para escribir
			
				registers[A3] <= WD3; // WD3 contiene el valor del registro 
			
			end
			
			registers[15] <= R15; // cambiar esto
			
		end
	
	end
	
	// lectura se hace en flanco negativo
	always_ff @(negedge clk or posedge rst) begin
	//always_ff @(*) begin
	
		if (rst) begin
		 // Reset behavior
			RD1_temp <= 16'h0;
			RD2_temp <= 16'h0;
			
		end 
		
		else begin
			RD1_temp <= registers[A1];
			RD2_temp <= registers[A2];
		end
	
	end
	
	assign RD1 = RD1_temp;
	assign RD2 = RD2_temp;

endmodule