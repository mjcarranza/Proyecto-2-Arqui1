module videoGen(
	input logic [9:0] x, y,
	output logic [7:0] r, g, b
);

	
	always @* begin
		{r, g, b} = {8'hFF, 8'h00, 8'h00};
	end
	
endmodule